module prueba(cornudo, raul);

input cornudo;
output raul;

endmodule