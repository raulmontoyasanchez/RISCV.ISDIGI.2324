module ALU_CONTROL(ALUOP, INSTRUCCION, ALUSELECT);
input [2:0]ALUOP;
input [3:0] INSTRUCCION;
output reg [3:0]ALUSELECT;

always @(ALUOP or INSTRUCCION)
if (ALUOP==2'b00)//RFORMAT
	begin
	case(INSTRUCCION)
	4'b0000: ALUSELECT=	4'b0000;//ADD
	4'b0001: ALUSELECT= 4'b0011; //DESPLAZAMIENTO IZQD
	4'b0010: ALUSELECT= 4'b0100; // MENOR QUE
	//4'b0011: ALUSELECT= 4'b????; // MENOR QUE UNSIGNED
	4'b0100: ALUSELECT= 4'b0111; // XOR
	4'b0101: ALUSELECT= 4'b0101; // DESPLAZAMIENTO DRCH
	4'b0110: ALUSELECT= 4'b0010; // OR
	4'b0111: ALUSELECT= 4'b0001; // AND
	4'b1000: ALUSELECT= 4'b0110;
	default: ALUSELECT = 4'b0000;
	endcase// SUB
	end
else if (ALUOP==2'b01)// RESTA(COMPARACION)
	 ALUSELECT = 4'b0110;
else if (ALUOP==2'b10)//SUMA(Direcciona memoria)
	 ALUSELECT= 4'b0000;
else
	ALUSELECT = 4'b0000;
	 

endmodule  

