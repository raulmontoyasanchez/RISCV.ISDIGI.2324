`timescale 1 ns/ 1 ps
module SINGLECYCLE();
logic CLK,RST;


TOP TOP_inst


endmodule