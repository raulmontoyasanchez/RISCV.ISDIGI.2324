module ALU_CONTROL();
input [1:0]ALUOP;
input [3:0] INSTRUCCION;
output reg [3:0]ALUSELECT;

always @(ALUOP or INSTRUCCION)
if (ALUOP=2'b00)//RFORMAT
	case(INSTRUCCION)
	4'b0000: ALUSELECT=	4'b0000;//SUMA
	4'b0001: ALU_SELECT= 4'b0001; //RESTA
else if (ALUOP=2'b01)//IFORMAT
	ALUSELECT = 4'b0001; //RESTA
else
	ALUSELECT==2'b00 
endmodule 