//MODULO DEL HAZARD DETECTION UNIT PARA EL CONTROL DE RIESGOS DEL DISEÑO PIPELINE DEL CORE

module HAZARD_DETECTION_UNIT(RS1_HDU, RS2_HDU, RD_EX, MEMREAD_EX, MUX_CONTROL_SELECT, REG_IF_ID_WRITE, PCWRITE);

//DECLARACION DE VARIABLES

//EX == PERTENECIENTE A ETAPA DE EJECUCION
//HDU == HAZARD DETECTION UNIT

input [4:0] RS1_HDU, RS2_HDU, RD_EX;
input MEMREAD_EX;

output MUX_CONTROL_SELECT, REG_IF_ID_WRITE, PCWRITE;

//CODIGO:

if (MEMREAD_EX && (RD_EX==RS1_HDU) or (RD_EX==RS1_HDU)
begin
	begin
	MUX_CONTROL_SELECT <= 1'b0;
	REG_IF_ID_WRITE <= 1'b0;
	PCWRITE <= 1'b0;
	end
else
	begin
	MUX_CONTROL_SELECT <= 1'b1;
	REG_IF_ID_WRITE <= 1'b1;
	PCWRITE <= 1'b1;
	end
end

endmodule 