module RAM (CLK, RESET_N, WRITE, READ, DATA_IN, ADDRESS, DATA_OUT);

//PARAMETROS

parameter TAM_POSICIONES=1024, TAM_PALABRA=32;	
//TAM_POSICIONES = N POSICIONES DE LA MEMORIA ; TAM_PALABRA = TAMANYO DE CADA POSICION DE MEMORIA
//DECLARACION DE VARIABLES


input CLK, RESET_N, WRITE, READ;
input [TAM_PALABRA-1:0] DATA_IN;
input [$clog2(TAM_POSICIONES)-1:0] ADDRESS;
output [TAM_PALABRA-1:0] DATA_OUT;

//MEMORIA RAM


reg [TAM_PALABRA-1:0]  [TAM_POSICIONES-1:0] MRAM;

//reg [TAM_PALABRA-1:0] DATA_OUT_AUX;

//CODIGO:

//LECTURA
assign DATA_OUT = (READ == 1'b1) ? MRAM[ADDRESS]  : 8'b0;

// ESCRITURA 
// ESCRIBIR : CUANDO WR = 1
 
always @(posedge CLK or negedge RESET_N)
 begin
	if (!RESET_N)
		MRAM <= '0;
		
	else if (WRITE) 
		MRAM[ADDRESS] <= DATA_IN;
			
 end
 
endmodule 