module TOP #(parameter ROM_INS=32, RAM_DATA=32, ROM_ADD=10, RAM_ADD=10) (CLK, RST);

//VARIABLES GENERALES
input CLK, RST;

//CABLES ROM
wire [ROM_ADD-1:0] ROM_ADDRESS;
wire [ROM_INS-1:0] ROM_INSTRUCTION;
//wire ROM_ENABLE;

//CABLES RAM
wire [RAM_DATA-1:0] RAM_DATAOUT;
wire [RAM_DATA-1:0] RAM_DATAIN;
wire [ROM_ADD-1:0] RAM_ADDRESS;
wire RAM_OUTPUT_ENABLE;
wire RAM_ENABLE_WR;

//RAM INSTANCIA
RAM RAM_INST(
.CLK(CLK),
.RSTa(RST),
.WR(RAM_ENABLE_WR), 
.OE(RAM_OUTPUT_ENABLE), 
.DATA_IN(RAM_DATAIN), 
.ADDRESS(RAM_ADDRESS), 
.DATA_OUT(RAM_DATAOUT)
);

//ROM INSTANCIA
ROM ROM_INST(
.READ_EN(1'b1),
.INS_ADDRESS(ROM_ADDRESS),
.INSTRUCTION_OUT(ROM_INTRUCTION)
);

//CORE INSTANCIA
CORE CORE_INST(
.CLK(CLK),
.RST_n(RST),
.DATA_IMEM(ROM_INTRUCTION),
.DATA_READ_DMEM(RAM_DATAOUT),
.DIR_IMEM(ROM_ADDRESS),
.DIR_DMEM(RAM_ADDRESS),
.DATA_WRITE_DMEM(RAM_DATAIN),
.READ(RAM_OUTPUT_ENABLE),
.WRITE(RAM_ENABLE_WR)
);

endmodule 