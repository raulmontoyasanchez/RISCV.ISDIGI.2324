module TOP (CLK, RESET_N, RAM_DATAOUT, RAM_DATAIN, RAM_ADDRESS);
//VARIABLES GENERALES
input CLK, RESET_N;

//CABLES ROM
wire [31:0] ROM_ADDRESS;
wire [31:0] ROM_INSTRUCTION;
wire READ, WRITE;
//wire ROM_ENABLE;

//CABLES RAM 
output wire [31:0] RAM_DATAOUT;
output wire [31:0] RAM_DATAIN;
output wire [31:0] RAM_ADDRESS;


//RAM INSTANCIA


RAM RAM_INST(
		.CLK(CLK),
		.RESET_N(RESET_N),
		.WRITE(WRITE), 
		.READ(READ),
		.DATA_IN(RAM_DATAIN),
		.DATA_OUT(RAM_DATAOUT),
		.ADDRESS(RAM_ADDRESS[11:2])

);

//ROM INSTANCIA
ROM ROM_INST(
.INS_ADDRESS(ROM_ADDRESS[11:2]),
.INSTRUCTION_OUT(ROM_INSTRUCTION),
.READ_EN(1'b1)
);

//CORE INSTANCIA
CORE CORE_INST(
.CLK(CLK),
.RESET_N(RESET_N),
.DATA_IMEM(ROM_INSTRUCTION),
.DATA_READ_DMEM(RAM_DATAOUT),
.DIR_IMEM(ROM_ADDRESS),
.DIR_DMEM(RAM_ADDRESS),
.DATA_WRITE_DMEM(RAM_DATAIN),
.READ(READ),
.WRITE(WRITE)
);

endmodule 