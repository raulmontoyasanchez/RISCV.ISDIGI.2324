module jajsjsjsdcbsxak


endmodule 